module not_14(
a,f
    );
    input wire [3:0]a;
    output wire [3:0]f;
    assign f = ~a ;
endmodule