/* Or gate with 2 1 bit inputs
Sum = a or b*/   /* */  //is used for multiline commmenting

module myor(a,b,y);

input a ,b;

output y;

assign y= a | b;

endmodule
//things in red mean preassigned things!!!