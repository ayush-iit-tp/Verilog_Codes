/* Or gate with 2 1 bit inputs
Sum = a or b*/   /* */  //is used for multiline commmenting

module mynot(a,y);

input a;

output y;

assign y= ~a;

endmodule
//things in red mean preassigned things!!!